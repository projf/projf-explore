// Project F: FPGA Graphics - Colour Test (Verilator SDL)
// (C)2022 Will Green, open source hardware released under the MIT License
// Learn more at https://projectf.io/posts/fpga-graphics/

`default_nettype none
`timescale 1ns / 1ps

module top_colour #(parameter CORDW=10) (  // coordinate width
    input  wire logic clk_pix,             // pixel clock
    input  wire logic sim_rst,             // sim reset
    output      logic [CORDW-1:0] sdl_sx,  // horizontal SDL position
    output      logic [CORDW-1:0] sdl_sy,  // vertical SDL position
    output      logic sdl_de,              // data enable (low in blanking interval)
    output      logic [7:0] sdl_r,         // 8-bit red
    output      logic [7:0] sdl_g,         // 8-bit green
    output      logic [7:0] sdl_b          // 8-bit blue
    );

    // display sync signals and coordinates
    logic [CORDW-1:0] sx, sy;
    logic de;
    simple_480p display_inst (
        .clk_pix,
        .rst_pix(sim_rst),
        .sx,
        .sy,
        /* verilator lint_off PINCONNECTEMPTY */
        .hsync(),
        .vsync(),
        /* verilator lint_on PINCONNECTEMPTY */
        .de
    );

    // screen dimensions (must match display_inst)
    localparam H_RES = 640;  // horizontal screen resolution
    localparam V_RES = 480;  // vertical screen resolution

    // determine colour from screen position
    logic [3:0] paint_r, paint_g, paint_b;
    always_comb begin
        if (sx < 256 && sy < 256) begin  // colour square in top-left 256x256 pixels
            paint_r = sx[7:4];  // 16 horizontal pixels of each red level
            paint_g = sy[7:4];  // 16 vertical pixels of each green level
            paint_b = 4'h4;     // constant blue level
        end else if (sx < H_RES-1 && sy < V_RES-1) begin  // otherwise dark blue
            paint_r = 4'h0;
            paint_g = 4'h1;
            paint_b = 4'h2;
        end else begin  // black in blanking interval
            paint_r = 4'h0;
            paint_g = 4'h0;
            paint_b = 4'h0;
        end
    end

    // SDL output (8 bits per colour channel)
    always_ff @(posedge clk_pix) begin
        sdl_sx <= sx;
        sdl_sy <= sy;
        sdl_de <= de;
        sdl_r <= {2{paint_r}};  // double signal width from 4 to 8 bits
        sdl_g <= {2{paint_g}};
        sdl_b <= {2{paint_b}};
    end
endmodule
